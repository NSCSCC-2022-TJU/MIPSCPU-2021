`include "defines.v"

module exe_stage (
    input  wire 					cpu_clk_50M,//闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺屻倝宕崟顐熷亾婵犳凹鏁嗛柡灞诲劚缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈敓锟�
    input  wire 					cpu_rst_n,
    // 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戞俊鐑芥晜閽樺澶勯梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁婀遍崗姗€寮ㄦ潏銊ヮ嚤闁跨噦鎷�
    // input   wire [`ALUTYPE_BUS	] 	exe_alutype_i,
    input   wire [`ALUOP_BUS	] 	exe_aluop_i,
    input   wire [`REG_BUS 		] 	exe_src1_i,
    input   wire [`REG_BUS 		] 	exe_src2_i,
    input   wire [`REG_ADDR_BUS ] 	exe_wa_i,
    input   wire 					exe_wreg_i,
    input	wire	                exe_mreg_i,
    input	wire [`REG_BUS	]	    exe_din_i,
    input	wire	                exe_whilo_i,
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垳绱掔€Ｑ冩櫛LO闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖娣灪缂嶅洭鏌ｉ幇闈涘妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁诡喗濞婇、鏇㈡晜閼恒儲顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼紒妯绘闂佽法鍣﹂幏锟�
    input	wire [`REG_BUS	]	    hi_i,
    input	wire [`REG_BUS	]	    lo_i,
    //闂傚倷娴囧▔鏇㈠窗閹邦喗鏆滈悗闈涙啞婵ジ鏌ら幇浣哥仭鐟滄妸鍥ㄧ厵濡炲楠搁崢鎾煛娴ｅ搫鏋戦柟宄版噹椤撳吋寰勭€ｎ偅顏熷┑掳鍊栭〃澶愬Υ閳ь剚淇婇幓鎺戭伃妤犵偛绻橀幃婊堟嚍閵夛附顏熺紓鍌欐祰鐏忔瑩宕滄ィ鍐┾拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箳缁岸寮伴敓锟�(add)
    input   wire                    mem2exe_whilo,
    input   wire [`DOUBLE_REG_BUS]  mem2exe_hilo,
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垳鈧懓瀚姗€寮查幖浣光拺閻犳亽鍔岄弸鎴︽煕閳轰焦鍤囨慨濠傘偢閹虫粌鈻撻崹顔芥澑濠电偞娼欓崥瀣偡閿旈敮鍋撳顒傜Ш鐎规洩缍佸浠嬵敇閻斿憡顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橀硸鍔廼闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垳绱掔仦鐐枔(add)
    input   wire                    wb2exe_whilo,
    input   wire [`DOUBLE_REG_BUS]  wb2exe_hilo,
    input   wire [`INST_ADDR_BUS ]  ret_addr,
    //闂傚倷娴囧▔鏇㈠窗鎼淬劍鍎戦柛鎾楀嫭娈伴梺褰掓？閻掞箓寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佽壘缂嶅﹪寮婚妸鈺傚亞闁稿本绋戦锟�
    input   wire [`REG_ADDR_BUS ] 	cp0_addr_i,
    input   wire [`REG_BUS ] 	    cp0_data_i,
    input   wire                    mem2exe_cp0_we,
    input   wire [`REG_ADDR_BUS ] 	mem2exe_cp0_wa,
    input   wire [`REG_BUS ] 	    mem2exe_cp0_wd,
    input   wire                    wb2exe_cp0_we,
    input   wire [`REG_ADDR_BUS ] 	wb2exe_cp0_wa,
    input   wire [`REG_BUS ] 	    wb2exe_cp0_wd,
    input   wire [`INST_ADDR_BUS ]  exe_pc_i,
    input   wire                    exe_in_delay_i,
    input   wire [`EXC_CODE_BUS ]   exe_exccode_i,

    // 闂備礁婀遍悷鎶藉炊閵婏附顏熼梻浣告啞閻燁垶宕戞繝鍋界喐鎷呴悜妯侯€涢柣鐔哥懃鐎氼剟顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐎涙绉堕梺鍛婂姈鐎笛呪偓姘炬嫹
    output  wire [`ALUOP_BUS] 	    exe_aluop_o,
    output  wire [`REG_ADDR_BUS] 	exe_wa_o,
    output  wire 					exe_wreg_o,
    output  wire [`REG_BUS]  	    exe_wd_o,
    output  wire	                exe_mreg_o,
    output	wire [`REG_BUS]	        exe_din_o,
    output	wire	                exe_whilo_o,
    output	wire [`DOUBLE_REG_BUS]	exe_hilo_o,
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш鐎规洘绮岄鍏煎緞鐎ｎ偅顏熼梻浣虹帛閻熻京妲愰弴鈧偓鍌烆敋閳ь剟鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣烘嚀閸ゆ牠骞忛敓锟�
    output wire                     exe2id_wreg,
    output wire [`REG_ADDR_BUS ]    exe2id_wa,
    output wire [`REG_BUS      ]    exe2id_wd,
    output wire                     exe2id_mreg,    
    //闂備礁婀遍悷鎶藉炊閵婏附顏熼梻浣告啞閻燁垶宕戞繝鍋界喐鎷呯化鏇熺亖闂傚倸鐗婄粙鎴濃枔閳哄懏鐓欏瀣閸樻挳鏌℃担瑙勫磳鐎殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉虹€规洘鍨甸オ浼村醇閻斿憡顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備胶鎳撻崵鏍箯閿燂拷
    output	wire	                stallreq_exe,
    //闂傚倷娴囧▔鏇㈠窗鎼淬劍鍎戦柛鎾楀嫭娈伴梺褰掓？閻掞箓寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佽壘缂嶅﹪寮婚妸鈺傚亞闁稿本绋戦锟�
    // output	wire	                cp0_re_o,
    output  wire [`REG_ADDR_BUS ] 	cp0_raddr_o,
    output	wire	                cp0_we_o,
    output  wire [`REG_ADDR_BUS ] 	cp0_waddr_o,
    output	wire [`REG_BUS]	        cp0_wdata_o,
    output  wire [`INST_ADDR_BUS ]  exe_pc_o,
    output	wire	                exe_in_delay_o,
    output  wire [`EXC_CODE_BUS ]   exe_exccode_o
    );

    // 闂備胶鍎甸弲婊堝箰閹惰棄鏋侀柟鎹愵嚙缁犳娊鏌曟径鍫濆鐟滄妸鍥ㄧ厵濡炲楠搁崢鎾煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煣濮橆剙鈧顢旈柆宥嗏拺閻犳亽鍔岄弸娑欎繆椤栨瑧顦﹂柍缁樻崌閹棄鈻撻幐搴㈩唶闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鐓欐い鎾卞妽鐎氾拷
    assign exe_aluop_o  =   exe_aluop_i;
    assign exe_mreg_o	=	exe_mreg_i;
    assign exe_din_o	=	exe_din_i;
    assign exe_whilo_o	=	exe_whilo_i;
    assign exe_pc_o     =   exe_pc_i;
    assign exe_in_delay_o=  exe_in_delay_i;
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш鐎规洘绮岄鍏煎緞鐎ｎ偅顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮樼偓瀚�
    assign exe2id_wreg = exe_wreg_i;
    assign exe2id_wa   = exe_wa_i;
    assign exe2id_mreg = exe_mreg_i;
    
    wire    [`REG_BUS ]         logicres;   //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏＄瑹椤栨瑧妫紓浣鸿檸閸欏啴寮ㄦ潏鈹惧亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閺佹捇鏁撻敓锟�
    wire	[`REG_BUS ]	        shiftres;   //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣告贡閺屽銆掗崷顓犵闁告稑鐡ㄩ悡銉╂煟閺傛寧鍟為柣蹇ｅ櫍閺岀喐顦版惔鈥冲箣闂佽桨鐒﹂幑鍥ь嚕椤掑嫬围闁糕剝顨忔导鎾绘⒒娴ｈ姤纭堕柛鐘冲姍瀵憡绻濆顒傤唵闂佽法鍣﹂幏锟�
    wire	[`REG_BUS ]	        moveres;    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ传閸曨厼闄嶉梺鑽ゅС濞村洭锝炴径灞稿亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備浇娉曢崳锕傚箯閿燂拷
    wire	[`REG_BUS ]	        hi_t;	    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧姀i闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖娣灪缂嶅洭鏌ｉ幇闈涘妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熺厱濠电姴绻戠€氾拷
    wire	[`REG_BUS ]	        lo_t;	    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧姌o闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖娣灪缂嶅洭鏌ｉ幇闈涘妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熺厱濠电姴绻戠€氾拷
    wire	[`REG_BUS ]	        arithres;	//闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш妤犵偛鐗撳鎾閳╁啯顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮樼偓瀚�
    wire	[`REG_BUS ]	        memres;	    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鎰佹綈缂佸锕畷濂稿Ψ閿旇姤顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鐓曠憸澶愬磻閿燂拷
    wire	[`REG_BUS ]	        cp0_t;      //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧妷p0闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖娣灪缂嶅洭鏌ｉ幇闈涘妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熺厱濠电姴绻戠€氾拷
    
    wire	[`DOUBLE_REG_BUS]	mulres;     //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш鐎殿喚鏁诲顕€宕奸悢鍛婎仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熺厵閺夊牄鍔嶇粈瀣煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱�(add)
    wire	[`DOUBLE_REG_BUS]	mulures;
    reg     [`DOUBLE_REG_BUS]   divres;      // 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш妤犵偛鐗撳鎾閳╁啯顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮樼偓瀚�

/*********************** 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш妤犵偞鍔欏畷鍫曨敆娴ｈ顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閿燂拷 begin*******************************/
    
    
    // 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈敓锟�
    wire                      signed_div_i;
    wire [`REG_BUS          ] div_opdata1;
    wire [`REG_BUS          ] div_opdata2;
    wire                      div_start;
    reg                       div_ready;

    assign stallreq_exe = 
                          (((exe_aluop_i == `MINIMIPS32_DIV) || (exe_aluop_i == `MINIMIPS32_DIVU))  && (div_ready == `DIV_NOT_READY))  ? `STOP : `NOSTOP;

    assign div_opdata1  = 
                          ((exe_aluop_i == `MINIMIPS32_DIV) || (exe_aluop_i == `MINIMIPS32_DIVU)) ? exe_src1_i : `ZERO_WORD;

    assign div_opdata2  = 
                          ((exe_aluop_i == `MINIMIPS32_DIV) || (exe_aluop_i == `MINIMIPS32_DIVU)) ? exe_src2_i : `ZERO_WORD;                                    
    assign div_start    = 
                          (((exe_aluop_i == `MINIMIPS32_DIV) || (exe_aluop_i == `MINIMIPS32_DIVU)) && (div_ready == `DIV_NOT_READY))  ? `DIV_START : `DIV_STOP; 

    assign signed_div_i = 
                          (exe_aluop_i == `MINIMIPS32_DIV ) ? 1'b1 : 1'b0; 

    wire   [34:0]                     div_temp;
    wire   [34:0]                     div_temp0;
    wire   [34:0]                     div_temp1;
    wire   [34:0]                     div_temp2;
    wire   [34:0]                     div_temp3;
    wire   [ 1:0]                     mul_cnt;

    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垳鈧懓瀚竟鍡欑矓閸ф鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備浇妗ㄩ悞锕傛偡閵夆晛鍚归柡宥庡幖缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囪尙顦柣鐘充航閸斿﹪鍩€椤掆偓椤戝鐛箛娑欏€婚柤鎭掑劜濞呫垽鏌ｉ悙瀵糕姇妞ゃ劍鍔楃槐鐐哄炊椤掆偓缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈敓锟�16闂備礁鎼崯顐︽偉婵傜ǹ鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛鏃戞Ч閹煎瓨绋愮划鐢告⒒娴ｈ姤纭堕柛鐘冲姍瀵憡绻濆顒傤唵闂佺粯鍨兼慨銈夊疾閹间焦鐓涘ù锝呮贡閹冲啴鏌涢妶鍡欏⒌妤犵偛绻橀幃婊堟嚍閵夛附顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備胶鎳撻崵鏍箯閿燂拷
    reg    [ 5:0]                     cnt;

    reg    [65:0]                     dividend;
    reg    [ 1:0]                     state;
    reg    [33:0]                     divisor;
    reg    [31:0]                     temp_op1;
    reg    [31:0]                     temp_op2;
    
    wire   [33:0]                     divisor_temp;
    wire   [33:0]                     divisor2;
    wire   [33:0]                     divisor3;
    
    assign divisor_temp = temp_op2;                   
    assign divisor2     = divisor_temp << 1;       //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熺厸闁割偆鍠愰ˉ鍫ユ煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕抽敃鍌氱闁跨噦鎷�
    assign divisor3     = divisor2 + divisor;      //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳鐐
    
    //dividend闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖杈剧到閺嬪牆顭跨捄渚剰妞ゅ骏鎷�32濠电偠鎻徊鐣岀矓瑜版帒鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳杈ㄥ殌妞ゎ厼娲らオ浼村醇閻斿憡顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箰閻ｏ繝骞嶉鐣岀Х闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠鸿櫣绛忛梺闈涚箞閸婃牠寮查幖浣哥骇闁绘劘鍩栫涵鑸点亜閿濆骸娅嶆鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閺屻劎鈧綆鍋掑Σ顖炴⒒娴ｈ姤纭堕柛鐘冲姍瀵憡绻濆顒傤唵缂備礁鑻绺眎dend[k:0]  
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш鐎殿喚鏁绘俊鎼佸煛閸屾稒顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉虹€规洖銈搁獮瀣晜閼恒儲顏熼梺鑽ゅ枑閻燂妇鏁幒鎾村劅婵犲﹤鐗嗙粻顖氼渻鐎ｎ亪顎楃紓鍌涘哺濮婅櫣鎹勯妸銉︾€鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒佽础濞寸媴绠撻獮瀣晜閼恒儲顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼捄铏圭瓘濠电偛鐬奸幉娌琩end[32:k+1]闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш鐎殿喚鏁绘俊鎼佸煛閸屾稒顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮樿鲸鍤€妞ゎ厼娲らオ浼村醇閻斿憡顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鍋ｉ悗锝冨妼閻忔煡鏌℃担瑙勫磳闁诡垰鐭傞、鏇㈡晬閸曨亣顩梻浣哥秺椤ユ捇寮绘径鎰？濠电姴娲﹂悡銉╂煟閺傛寧鍟為柣蹇ｅ櫍閺岀喐顦版惔鈥冲箣闂佽桨鐒﹂幑鍥ь嚕椤掑嫬围闁糕剝顨忔导鎾绘⒒娴ｈ姤纭堕柛鐘冲姍瀵憡绻濆顒傤唵闂佺粯鍨兼慨銈夊疾閹间焦鐓ラ柣鏇炲€圭€氾拷  
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏㈢矙鐠恒劊鍋ｉ梻浣瑰缁诲倻鎹㈤幋鐘亾濮橀硸鍔奿vidend闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘32濠电偠鎻徊鐣岀矓瑜版帒鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繗鍩栭幈銊╂晲閸涱垳顔掗梺杞扮劍閹歌顭囬鍡樺磯妞ゎ厽鍨跺▓浼存⒑瑜版帩妫戦柛蹇旓耿瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鐓涢柛鎰╁妿閸╋綁鏌℃担瑙勫鞍缂佹鍠栨俊鐑芥晝閳ь剟寮ィ鍐╃厵濡炲楠搁崢鎾煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煥閻曞倹瀚�
    assign div_temp0 = {1'b000,dividend[63:32]} - {1'b000,`ZERO_WORD};  //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸娆愩亜閺囩姴啸闁诡噮鍣ｉ、鏇㈡晜閼恒儲顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閿燂拷 0 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻缂佹ɑ娅㈤梺璺ㄥ櫐閹凤拷
    assign div_temp1 = {1'b000,dividend[63:32]} - {1'b0,divisor};       //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸娆愩亜閺囩姴啸闁诡噮鍣ｉ、鏇㈡晜閼恒儲顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閿燂拷 1 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻缂佹ɑ娅㈤梺璺ㄥ櫐閹凤拷
    assign div_temp2 = {1'b000,dividend[63:32]} - {1'b0,divisor2};      //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸娆愩亜閺囩姴啸闁诡噮鍣ｉ、鏇㈡晜閼恒儲顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閿燂拷 2 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻缂佹ɑ娅㈤梺璺ㄥ櫐閹凤拷
    assign div_temp3 = {1'b000,dividend[63:32]} - {1'b0,divisor3};      //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸娆愩亜閺囩姴啸闁诡噮鍣ｉ、鏇㈡晜閼恒儲顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閿燂拷 3 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻缂佹ɑ娅㈤梺璺ㄥ櫐閹凤拷
    
    assign div_temp  = (div_temp3[34] == 1'b0 ) ? div_temp3 : 
                       (div_temp2[34] == 1'b0 ) ? div_temp2 : div_temp1;
                      
    assign mul_cnt   = (div_temp3[34] == 1'b0 ) ? 2'b11 : 
                       (div_temp2[34] == 1'b0 ) ? 2'b10 : 2'b01;
    
    always @ (posedge cpu_clk_50M) begin
        if (cpu_rst_n == `RST_ENABLE) begin
            state         <= `DIV_FREE;
            div_ready     <= `DIV_NOT_READY;
            divres       <= {`ZERO_WORD,`ZERO_WORD};
        end else begin
        case (state)
    //*******************   DIV_FREE闂備胶绮灙闁糕晜鐗犻崺鈧い鎺戯攻鐎氾拷    ***********************  
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備浇娉曢崳锕傚箯閿燂拷  
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘1闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鎰佹綈闁逛究鍔庨埀顒婄秵閸犳寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佽壘缂嶅﹪寮婚妸鈺傚亜闁告稑锕︽导鍕⒑瑜版帩妫戦柛蹇旓耿瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬪孩銇勯锝嗙闁轰礁绉撮悾婵嬪礋椤掍焦顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫瑥鈹戦悙鍙夊枠闁轰焦鎹囬弫鎾绘晸閿燂拷0闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鎰佹綈缂佸锕畷濂稿Ψ閿旇姤顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾瑰姽ivByZero闂備胶绮灙闁糕晜鐗犻崺鈧い鎺戯攻鐎氾拷  
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘2闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鎰佹綈闁逛究鍔庨埀顒婄秵閸犳寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佽壘缂嶅﹪寮婚妸鈺傚亜闁告稑锕︽导鍕⒑瑜版帩妫戦柛蹇旓耿瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬪孩銇勯锝嗙闁轰礁绉撮悾婵嬪礋椤掍焦顏熼梻浣筋潐濡炲潡宕㈡ィ鍐炬晢闁哄被鍎辩粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁婀遍弻澶娿€掗崷顓熷闁跨噦鎷�0闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鎰佹綈缂佸锕畷濂稿Ψ閿旇姤顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾瑰姽ivOn闂備胶绮灙闁糕晜鐗犻崺鈧い鎴ｆ硶缁愭棃鏌℃担瑙勫磳鐎殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖溾偓鐟板閸嬪﹤顭囧Δ鍛拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箳缁碍鍒婂娑欑箾閹寸偞鎯堥柟鍑ゆ嫹0闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鐐  
    //     闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏犵暋閺夎法绱﹂梻浣告啞閸垶宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垻鎷犻幓鎺濇缂傚倷鐒︾粙鏍綖婢跺备鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴犳喐闁箑娅嶆鐐差槺閳ь剨缍嗛崑鍕敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻閸撲礁宕ュ銈嗘尵婵參宕濆⿰鍫熺厵濡炲楠搁崢鎾煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹀┑鐐村灦閹歌顪冩禒瀣瀬闁规崘顕уΛ姗€鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳鎰佹綈缂佸锕畷濂稿Ψ閿旇姤顏熼梻浣圭湽閸斿苯螞濞嗘挸鑸瑰┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鏃€銇勮箛锝勭敖缂侇喚鏁搁幉鎾礋椤愵偂绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬪秹鏌ら悡搴㈡崳闁归濮鹃ˇ鎶芥倵濮橆剛绉洪柡灞诲姂閹垹煤鐠囧弶顓婚梻渚€娼уΛ鎾箯閿燂拷  
    //     闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻缂佹ê娈熼梺闈涱槶閸庨亶鎮℃穱顦弙isor闂傚倷娴囧▔鏇㈠窗鎼淬們浜归柕濞炬櫆閺呮煡鐓崶銊︾叆妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏㈡嫚濞村鐎煎┑鐐存綑閸氬鎮烽敂閿亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備胶鎳撻崲鏌ュ床閺屻儲绠掔紓鍌欑瀵爼鏌ч崐淇癲end闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖杈剧到閺嬪牆顭跨捄渚剰妞ゅ骏鎷�32濠电偠鎻徊鐣岀矓瑜版帒鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ骏鎷�  
    //     闂備礁鎲￠崹闈浳涘┑瀣瀬闁规崘顕уΛ姗€鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崨濠勬噽闁稿妫濋妴鍌烆敋閳ь剟鐛箛娑欐啣闁稿本绮犳导鍥⒒娴ｈ姤纭堕柛鐘虫礃缁绘盯宕堕埡浣圭€虫繝銏ｆ硾椤戝懘顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閺佹捇鏁撻敓锟�  
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘3闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶姊洪崹顕呭剳婵﹪绠栧铏规崉閵娿儲鐎婚悷婊嗗焽閸旀垵顕ｉ鍕ч柛鈩冾殢娴兼捇姊绘担鑺ョ《闁哥姴姘﹂妵鎰板Ω瑜忔す鎶芥偡濞嗗繐顏╂い蹇撶埣濮婅櫣鎹勯妸銉︾€鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏＄附婢跺绋愰梻浣瑰缁嬫垿鎯岄崒鐐叉瀬闁规崘顕уΛ姗€鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛鏇犵煔閻庡厜鏆ready濠电偞鍨堕幖顐﹀箯閿燂拷0闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垳绱掔仦绛嬪悪vres濠电偞鍨堕幖顐﹀箯閿燂拷0  
    //*********************************************************** 
              `DIV_FREE: begin                       //DIV_FREE
                  if(div_start == `DIV_START) begin
                      if(div_opdata2 == `ZERO_WORD) begin        // 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鎰佹綈缂佸顦甸弫鎾绘晸閿燂拷0
                          state <= `DIV_BY_ZERO;
                      end else begin                            // 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鎰佹綈缂佸顦甸弫鎾绘晸閿燂拷0
                          state <= `DIV_ON;
                          cnt   <= 6'b000000;
                        
                        if(exe_aluop_i == `MINIMIPS32_DIV) begin
                            if(div_opdata1[31] == 1'b1 ) begin
                                temp_op1 = ~div_opdata1 + 1;    // 闂備礁鎲￠悷锕傛偋閻樿鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垺绻涢幘鏉戞惛闁稿孩鎸抽、姘堪閸繄顔嗛梺缁樺灱婵倝寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佺啲閹凤拷
                            end else begin
                                temp_op1 = div_opdata1;
                            end
                            if(div_opdata2[31] == 1'b1 ) begin
                                temp_op2 = ~div_opdata2 + 1;    // 闂備礁鎲￠悷锕傛偋閻樿鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垺绻涢幘鏉戞惛闁稿孩鎸抽、姘堪閸繄顔嗛梺缁樺灱婵倝寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佺啲閹凤拷
                            end else begin
                                temp_op2 = div_opdata2;
                            end
                        end

                        else begin//(exe_aluop_i == `MINIMIPS32_DIVU)
                            temp_op1 = div_opdata1;
                            temp_op2 = div_opdata2;
                        end
                        
                        dividend        <= {`ZERO_WORD,`ZERO_WORD};
                        dividend[31:0]  <= temp_op1;
                        divisor         <= temp_op2;
                    end
                end else begin     // 婵犵數鍋涢惌澶屾崲濠靛鏋侀柟鎹愵嚙閻銇勯幇鈺佺仼闁活煉绻濋弻鐔风暋閺夋寧些濡炪値鍋呴崝娆撳蓟閵娾晜鍋勯柛娑橈功娴煎嫰姊鸿ぐ鎺濇闁稿繑锕㈠顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳鐐
                        div_ready  <= `DIV_NOT_READY;
                        divres <= {`ZERO_WORD,`ZERO_WORD};
                end              
              end

    //*******************   DivByZero闂備胶绮灙闁糕晜鐗犻崺鈧い鎺戯攻鐎氾拷    ********************  
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻閼告娼熺紓渚囧亞閹规墪yZero闂備胶绮灙闁糕晜鐗犻崺鈧い鎴ｆ硶缁愭棃鏌℃担瑙勫磳鐎殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煣濮橆剙鈧鎮块崟顖涚厽闁冲搫鍊圭亸锕傛煛娴ｈ宕屾鐐村浮婵＄兘鏁傞悾灞肩磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂缁傛vEnd闂備胶绮灙闁糕晜鐗犻崺鈧い鎴ｆ硶缁愭棃鏌℃担瑙勫磳鐎殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備浇顫夊鍧楀储娴犲鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐瀵爼鎮欓幓鎺旀闂佺懓鍤栭幏锟�0  
    //*********************************************************** 
              `DIV_BY_ZERO: begin               //DivByZero
                 dividend <= {`ZERO_WORD,`ZERO_WORD};
                  state    <= `DIV_END;                 
              end

    //*******************   DivOn闂備胶绮灙闁糕晜鐗犻崺鈧い鎺戯攻鐎氾拷      ***********************  
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘1闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゆ惞鐠団剝鐐妌t闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌у顒€鈧晫绮堥敓锟�16闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鎰佹綈缂佸锕畷濂稿Ψ閿旇姤顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剚璐＄紒顔肩墕鐓ゆい蹇撴噺濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲啰鏆氶梻浣告啞閸垶宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁婀遍崗姗€寮ㄩ柆宥嗗剦闁告稑鐡ㄩ悡銉╂煟閺傚灝妲荤€点倖妞介弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閺屻劎鈧綆鍋掑Σ锟�  
    //    闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箳缁氨鈧厜鏆temp濠电偞鍨堕幐璇差渻娴犲鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳鎰佹綈缂佸锕畷濂稿Ψ閿旇姤顏熼梻浣告啞閹歌崵鈧瑳鍥舵晝闁兼祴鏅涢弸鍫濐熆鐠轰警鍎忔い蹇撶埣濮婅櫣鎹勯妸銉︾€鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻缂佹ɑ娅㈤梺璺ㄥ櫐閹凤拷0闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鐐  
    //    闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鏃傜磼閸屾凹鍚檝_temp濠电偞鍨堕幐璇差渻娴犲鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳鎰佹綈缂佸锕畷濂稿Ψ閿旇姤顏熼梻浣告啞閹歌崵鈧瑳鍥舵晝闁兼祴鏅涢弸鍫濐熆鐠轰警鍎忔い蹇撶埣濮婅櫣鎹勯妸銉︾€鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻缂佹ɑ娅㈤梺璺ㄥ櫐閹凤拷1闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垳绱掔仦绛嬪悪vidend  
    //    闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏㈡嫚濞村鐎煎┑鐐存綑閸氬鎮烽敂閿亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼紒妯哄壒濡炪倖鍔戦崹褰掓儍閿熺姵鐓欏瀣閻掑潡鏌℃担鍓插剶闁诡啫鍥ㄦ櫢闁绘ǹ娅曞▍銏ゆ⒑閸濆嫬鈧爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箰閻ｏ繝鎮ч崼婵冨亾闁秵鐓涢柛鎰╁妿閸╋綁鏌℃担瑙勫磳鐎殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖滅磼鐎ｅ灚顫梫On闂備胶绮灙闁糕晜鐗犻崺鈧い鎴ｆ硶缁愭棃鏌℃担瑙勫磳鐎殿噮鍓熸俊鍫曞幢濡ゅ﹣绱nt闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘1闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘  
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘2闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゆ惞鐠団剝鐐妌t濠电偞鍨堕幖顐﹀箯閿燂拷16闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鎰佹綈缂佸锕畷濂稿Ψ閿旇姤顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剚璐＄紒顔肩墕鐓ゆい蹇撴噺濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲啰鏆氶梻浣告啞閸垶宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熺叆婵犲﹤鍟扮粔娲煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕抽敃鍌氱闁跨噦鎷�  
    //    闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囪尙顔屽銈嗘尵閸犲酣寮ィ鍐╃厵濡炲楠搁崢鎾煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂鐠鸿　妲堥柟缁㈠灠娴滈箖姊绘担鑺ョ《闁哥姵鍔欏鍛婄節濮橆剛顔嗛梺鐐壘閸婂顢旈柆宥嗏拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣告贡閺屽銆掗崷顓犱笉闁绘劗鍎ら悡銉╂煟閺傛寧鍟為柣蹇ｅ櫍閺岀喐顦版惔鈥冲箣闂佽桨鐒﹂幑鍥ь嚕椤掑嫬围闁糕剝顨忔导鎾绘⒒娴ｈ姤纭堕柛鐘冲姍瀵娊鍩€椤掑嫭鐓曢柟瀛樼懃閳ь剚鐗滈埀顒佽壘缂嶅﹪寮婚妸鈺傚亜闁诡垱婢橀婊堟⒑閸濆嫬鈧爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁诡啫鍥ㄥ亜闁稿繐鍚嬪▍銏ゆ⒑閸濆嫬鈧爼宕愰弽顐熷亾濮橆剛绉洪柟铏崌瀹曠喖妫冨☉妯锋寗闂備礁婀遍崗姗€藟閹捐埖鏆滈柛褎顨嗛悡銉╂煟閺傛寧鍟為柣蹇ｅ櫍閺岀喐顦版惔鈥冲箣闂佽桨鐒﹂幑鍥ь嚕椤掑嫬围闁糕剝顨忔导鎾绘⒑閻戔晜娅呯紒缁橈耿瀵偊骞樼紒妯绘闂佽法鍣﹂幏锟�  
    //    闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇寮绘径鎰瀭闁规儼濮ら悡銉╂煟閺傛寧鍟為柣蹇ｅ櫍閺岀喐顦版惔鈥冲箣闂佽桨鐒﹂幑鍥ь嚕椤掑嫬围闁糕剝顨忔导鎾绘⒑缂佹ü绶遍柛娆忓暣瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏㈢矙鐠恒劍鐎俊鐐€曠换鎰偓娑掓櫇閳ь剚鑹剧紞濠囧蓟閵娾晜鍋勯柛娑橈功娴煎嫰姊鸿ぐ鎺濇闁稿繑锕㈠顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箲椤︾増鎯旈埦鈧幏顐︽⒒娴ｈ姤纭堕柛鐘冲姍瀵憡绻濆顒傤唵闂備礁鐏濋鍡涘磿閸洘鐓ユ繝闈涙缁犳煡鎮楀顒傜Ш闁诡垯绶氶、鏇㈡晜閼恒儲顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼捄铏圭瓘濠电偛鐬奸幉娌琩end闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖杈剧到閺嬪牆顭跨捄渚剰妞ゅ骏鎷�32濠电偠鎻徊鐣岀矓瑜版帒鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳鐐  
    //    闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇銈惉姝穒dend闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖娣妽椤ュ牓鏌嶉崫鍕偓鎼侇敂閿燂拷32濠电偠鎻徊鐣岀矓瑜版帒鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖奸弻娑橆潩椤掍焦鎷卞┑锛勫仜閸婂潡寮婚妸鈺傚亜闁告稑锕︽导鍕⒑瑜版帩妫戦柛蹇旓耿瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂缁傛vEnd闂備胶绮灙闁糕晜鐗犻崺鈧い鎴ｆ硶缁愭棃鏌℃担瑙勫磳鐎殿噮鍓熸俊鍫曞幢濡ゅ﹣绱�  
    //***********************************************************
              `DIV_ON: begin               //DivOn
                  if(cnt != 6'b100010) begin    //cnt闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌у顒€鈧晫绮堥敓锟�16闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒佽础缂侇喖鐗嗙叅妞ゅ繐鎳忓▍銏ゆ⒑閸濆嫬鈧爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍐殮闂備礁鎲￠崹顖炲磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣告贡閸忔﹢寮ㄩ柆宥嗗剦闁告稑鐡ㄩ悡銉╂煟閺傚灝妲荤€点倖妞介弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備胶鎳撻崵鏍箯閿燂拷
                    if(div_temp[34] == 1'b1) begin
                        //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛憸缁辨帡宕ｆ径鎰儍v_temp[32]濠电偞鍨堕幖顐﹀箯閿燂拷1闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒佽础缂侇喖鐗嗙叅妞ゅ繐鎳忓▍銏ゆ⒑閸濆嫬鈧爼宕愰弽顐熷亾濮橀硸鍔歩nuend-n闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏犵暋閺夎法绱﹂梻浣哥枃濡嫰骞婅箛鏇楀亾濮橆剛绉洪柡灞诲姂閹倝宕掑☉姗嗕紦0闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘  
                          //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垳绱掔仦绛嬪悪vidend闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣告贡閺屽銆掗崷顓犲崥閻庢稒蓱婵鈧箍鍎遍ˇ浼村疾閹间焦鐓涢柛灞久埀顒佺墱閳ь剚鑹剧紞濠囧蓟閵娾晜鍋勯柛娑橈功娴煎嫰姊鸿ぐ鎺濇闁稿繑锕㈠顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸娑㈡煕濞嗘劖銇濈€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閼哥數绠剧€光偓鐎ｎ剛鐦堥梺杞扮劍閹瑰洤鐣烽敐澶樻晝闁靛鍠栧▓婵嬫⒑瑜版帩妫戦柛蹇旓耿瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銈夊磼濞戞﹩浼�  
                          //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐瀵爼鎮欑仦鍌欑钵缂備線纭搁崳锝夌嵁韫囨稒鍊婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳杈ㄥ殌妞ゎ偅绻堝畷锝嗗緞鐎ｎ兛绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囪尙顔屽銈嗘尰缁诲嫭绋夐弻銉︾厵濡炲瀛╅悞鍧楁煛娴ｅ壊鍎旈柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鍋ｉ悗锝庝憾閸庢棃鏌℃担瑙勫磳鐎殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉虹€殿喕绮欓弫鎾绘偐閾忣偅顏熼梻鍌欒兌婢ф顢欓弽顓炵？闂侇剙绉寸粻鐔兼倵閿濆骸浜滄い蹇撶埣濮婅櫣鎹勯妸銉︾彚闂佺懓鍤栭幏锟�0闂佸搫顦弲娆戝垝濞嗘挸鏋侀柟鎹愵嚙缁犳娊鏌曟竟顖氭湰濞堜即姊鸿ぐ鎺濇闁稿繑锕㈠顐﹀箻鐠囪尙鐓戝銈嗗姂閸婃垿鍩€椤掆偓椤戝鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳鐐
                        dividend <= {dividend[63:0] , 2'b00};
                    end else begin
                        //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛憸缁辨帡宕ｆ径鎰儍v_temp[32]濠电偞鍨堕幖顐﹀箯閿燂拷0闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒佽础缂侇喖鐗嗙叅妞ゅ繐鎳忓▍銏ゆ⒑閸濆嫬鈧爼宕愰弽顐熷亾濮橀硸鍔歩nuend-n闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熷仯闁搞儺鐓夐懓鍧楁煛娴ｈ宕岄柡浣规崌閺佹捇鏁撻敓锟�  
                          //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ㄩ悤鍌涘0闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸宥夋煠閻撳酣鍙勭€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴⒑閸噮鍎忛柡鍛櫅闇夐柛蹇氬亹閹冲嫰鎮楀顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鏃堟煟閹垮啫浜濋悗鐢靛帶閳诲酣骞囬澶夌处闂備胶鍘ч崢鏍濮樿泛鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐎涙ê顫℃繝銏ｆ硾閹芥粍绋夐弻銉︾厵濡炲楠搁崢鎾煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱︽繝娈垮枟閿氱€殿喖鐖煎鍛婄節濮橆剛顔嗛梺缁樺灱婵倝寮查幖浣圭叆闁绘洖鍊圭€氾拷  
                          //濠电偞鍨堕幐鎾磻閹剧粯鈷戦悹鎭掑妼閺嬫瑥鈹戦悙鍙夊窛闁哥姴锕ュ鍕偓锝庝憾娴兼捇姊绘担鑺ョ《闁哥姵鍔欏鍛婄節濮橆剛顔嗛梺缁樺灱婵倝寮茬粙瑁も偓鎺戭潩閵夈儱濮曢梺鍝ュ仜椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囪尙鐓戝銈嗗姦閸撴稓绮旈崼鏇熺厵鐎瑰嫭婢樺Σ濠氭煙椤旇姤宕岀€殿噮鍣ｅ畷濂稿即閻斿憡顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮樼偓瀚�1闂佸搫顦弲娆戝垝濞嗘挸鏋侀柟鎹愵嚙缁犳娊鏌曟竟顖氭湰濞堜即姊鸿ぐ鎺濇闁稿繑锕㈠顐﹀箻鐠囪尙鐓戝銈嗗姂閸婃垿鍩€椤掆偓椤戝鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳鐐 
                        dividend <= {div_temp[31:0] , dividend[31:0] , mul_cnt};
                    end
                    cnt <= cnt + 2;
                end else begin    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺屸剝鎷呴崷顓熷櫑闂佹悶鍊栭悧鐘荤嵁韫囨稒鍊婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣烘嚀閸ゆ牠骞忛敓锟�
                
                if(exe_aluop_i == `MINIMIPS32_DIV) begin
                    if((div_opdata1[31] ^ div_opdata2[31]) == 1'b1) begin
                        dividend[31:0] <= (~dividend[31:0] + 1);    // 闂備礁鎲￠悷锕傛偋閻樿鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垺绻涢幘鏉戞惛闁稿孩鎸抽、姘堪閸繄顔嗛梺缁樺灱婵倝寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佺啲閹凤拷
                    end
                    if((div_opdata1[31] ^ dividend[65]) == 1'b1) begin              
                        dividend[65:34] <= (~dividend[65:34] + 1);    // 闂備礁鎲￠悷锕傛偋閻樿鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垺绻涢幘鏉戞惛闁稿孩鎸抽、姘堪閸繄顔嗛梺缁樺灱婵倝寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佺啲閹凤拷
                    end
                end//`MINIMIPS32_DIV闂傚倷娴囧▔鏇㈠窗閹邦喗鍠嗛柨鏃傛櫕閳绘梻鈧箍鍎卞Λ娆撳汲椤撱垺鐓欓柟缁樺俯閸庢劙鎮楀槌栧妸ividend
                
                state <= `DIV_END;        //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧剾ivEnd闂備胶绮灙闁糕晜鐗犻崺鈧い鎺戯攻鐎氾拷 
                cnt   <= 6'b000000;       //cnt闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳鐐         
               end
              end

     //*******************   DivEnd闂備胶绮灙闁糕晜鐗犻崺鈧い鎺戯攻鐎氾拷    ***********************  
     //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゆ惞鐠団剝鎹秈vres闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖娣妼缁€宀勬煃閳轰礁鏆欐い蹇撶埣濮婅櫣鎹勯妸銉︾€鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳鐐64濠电偠鎻徊鐣岀矓瑜版帒鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊虹捄銊ユ珢闁瑰嚖鎷�32濠电偠鎻徊鐣岀矓瑜版帒鏋侀柟鍓х帛閸ゅ秹鏌曟径鍫濆姎濞存粌鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈敓锟�32濠电偠鎻徊鐣岀矓瑜版帒鏋侀柟鍓х帛閸ゅ秹鏌曟径鍫濆姎濞存粌鐖煎铏规崉閵娿儲鐎鹃梺鍝勬閸嬫捇姊洪幐搴ｇ畵缂佺粯鍨归埀顒佺啲閹凤拷  
     //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熺參婵☆垳绮粈瀣煛娴ｈ灏电€垫澘锕ら埢浠嬫偡閸椾拷eady濠电偞鍨堕幐楣冩儊濮濓箼ResultReady闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒佽础缂侇喖鐗嗙叅妞ゅ繐鎳忓▍銏ゆ⒑閸濆嫬鈧爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁诡喚鍋ゅ畷濂稿即閻斿憡顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉虹€规洩绻濋獮姗€顢欓懞銉︻仧缂傚倷娴囨禍顒勫磻閹稿簼绻嗘い鏍ュ€楃弧鈧梺杞扮劍閹瑰洤顕ｉ鍕ч柛鈩冾殢娴硷拷  
     //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧剾ivStop闂傚倷娴囧▔鏇㈠窗閺囥垹绀堝┑鍌溓归惌妤呮煕閹存瑥鈧绮旈崼鏇熺厵濡炲楠搁崢鎾煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱X婵犵妲呴崹鐣屾崲濠靛鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳槌栧剾ivStop闂傚倷娴囧▔鏇㈠窗閺囥垹绀堝┑鍌氭啞閸嬫牠鎮楀☉娅亪顢旈崼鏇熺厸闁告劑鍔庨崺锝夋煛娴ｈ宕岀€殿噮鍓熸俊鍫曞幢濡ゅ﹣绱IV婵犵妲呴崹鐣屾崲濠靛鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繗鍩栭幈銊ノ熺拠鎻掝潚闂佽桨鐒﹂幐鎯ｉ幇顔惧暗閻庢稓锕狥REE闂備胶绮灙闁糕晜鐗犻崺鈧い鎺戯攻鐎氾拷  
     //********************************************************** 
              `DIV_END: begin               //DivEnd
               divres <= {dividend[65:34], dividend[31:0]};  
               div_ready  <= `DIV_READY;
               if(div_start == `DIV_STOP) begin
                      state         <= `DIV_FREE;
                    div_ready     <= `DIV_NOT_READY;
                    divres      <= {`ZERO_WORD,`ZERO_WORD};
               end
              end
          endcase
        end
    end
/*********************** 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш妤犵偞鍔欏畷鍫曨敆娴ｈ顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閿燂拷 end*********************************/ 


    //闂傚倷娴囧▔鏇㈠窗鎼淬劍鍎戦柛鎾楀嫭娈伴梺褰掓？閻掞箓寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佽壘缂嶅﹪寮婚妸鈺傚亞闁稿本绋戦锟�
    assign cp0_we_o = 
        (exe_aluop_i==`MINIMIPS32_MTC0)?1'b1:1'b0;
    assign cp0_wdata_o = 
        (exe_aluop_i==`MINIMIPS32_MTC0)?exe_src2_i:`ZERO_WORD;
    assign cp0_waddr_o = cp0_addr_i;
    assign cp0_raddr_o = cp0_addr_i;
    // assign cp0_re_o = 
    //     (exe_aluop_i==`MINIMIPS32_MFC0)?1'b1:1'b0;
    //闂傚倷娴囧▔鏇㈠窗鎼淬們浜归柕濞у嫬顎涢柣鐔哥懃鐎氼剟顢旈崼鏇熲拺閻犳亽鍔岄弸娆愩亜椤愶綆娈滅€规洘鐟╂俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾汇偑閻拷0闂傚倷娴囧▔鏇㈠窗鎼淬們浜归柕濞р偓閸嬫捇妫冨☉姗嗕紓闂佽妞挎禍顏堢嵁韫囨稒鍊婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш鐎规洘顨婇崺鈧い鎺戝閻撱儵鏌ｉ弬鎸庡暈闁诲浚鍣ｉ弻鐔割槹鎼粹€冲箣闂佽桨鐒﹂幑鍥ь嚕椤掑嫬围闁糕剝顨忔导鎾绘⒒娴ｈ姤纭堕柛鐘冲姍瀵憡绻濆顒傤唵缂備礁鑻悰锟�0闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖娣灪缂嶅洭鏌ｉ幇闈涘妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熺厱濠电姴绻戠€氾拷
    assign cp0_t = //(cp0_re_o!=`READ_ENABLE)?`ZERO_WORD:
        (mem2exe_cp0_we==`WRITE_ENABLE && mem2exe_cp0_wa==cp0_raddr_o)?mem2exe_cp0_wd:
        (wb2exe_cp0_we==`WRITE_ENABLE && wb2exe_cp0_wa==cp0_raddr_o)?wb2exe_cp0_wd:cp0_data_i;

    
    // 闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧妴luop闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏＄瑹椤栨瑧妫紓浣鸿檸閸欏啴寮ㄦ潏鈹惧亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閿燂拷
    assign logicres = 
        (exe_aluop_i == `MINIMIPS32_AND ) ? (exe_src1_i & exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_ORI ) ? (exe_src1_i | exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_OR  ) ? (exe_src1_i | exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_NOR ) ? ~(exe_src1_i | exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_XOR ) ? (exe_src1_i ^ exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_ANDI) ? (exe_src1_i & exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_XORI) ? (exe_src1_i ^ exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_LUI ) ? exe_src2_i : `ZERO_WORD;
        
    
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧妴luop闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣告贡閺屽銆掗崷顓犵闁告稑鐡ㄩ悡銉╂煟閺傛寧鍟為柣蹇ｅ櫍閺岀喐顦版惔鈥冲箣闂佽桨鐒﹂幑鍥ь嚕椤掑嫬围闁糕剝顨忔导锟�
    assign shiftres = 
        (exe_aluop_i == `MINIMIPS32_SRL ) ? (exe_src2_i >> exe_src1_i):
        (exe_aluop_i == `MINIMIPS32_SRA ) ? $signed(($signed(exe_src2_i)) >>> exe_src1_i):
        (exe_aluop_i == `MINIMIPS32_SLLV) ? (exe_src2_i << exe_src1_i[4:0]):
        (exe_aluop_i == `MINIMIPS32_SRLV) ? (exe_src2_i >> exe_src1_i[4:0]):
        (exe_aluop_i == `MINIMIPS32_SRAV) ? $signed(($signed(exe_src2_i)) >>> exe_src1_i[4:0]):
        (exe_aluop_i == `MINIMIPS32_SLL ) ? (exe_src2_i << exe_src1_i) : `ZERO_WORD;
    
   //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧妴luop闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鏃堟倵濮橆厾銆掗柟宄邦儑閹叉挳宕熼顐＄处闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋綁顢樿娴滅偞銇勯敐搴℃珝妤犵偛绻橀幃婊堟嚍閵夛附顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕楅崗鐓庢珴缂備胶鍋撳姗€藝閹殿喒鍋撳槌栧劉ILO闂傚倷娴囧▔鏇㈠窗瀹ュ鍤戦幖娣灪缂嶅洭鏌ｉ幇闈涘妞ゅ繐鐖煎铏规崉閵娿儲鐎鹃梺鍝勵儏椤兘鐛箛娑欏€婚柤鎭掑劜濞呫垽姊洪崫鍕偓鍫曞磹閺嶎偀鍋撳顒傜Ш鐎规洘鍔欓弫鎾绘晸閿燂拷(MTHI,MTLO闂備礁婀辨灙婵炲樊鍙冨顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈敓锟�)
    assign hi_t =   
                    (mem2exe_whilo==`WRITE_ENABLE) ? mem2exe_hilo[63:32]:
                    (wb2exe_whilo==`WRITE_ENABLE) ? wb2exe_hilo[63:32] : hi_i;
    assign lo_t =   
                    (mem2exe_whilo==`WRITE_ENABLE) ? mem2exe_hilo[31:0]:
                    (wb2exe_whilo==`WRITE_ENABLE) ? wb2exe_hilo[31:0] : lo_i;

    assign moveres = 
        (exe_aluop_i == `MINIMIPS32_MFHI) ? hi_t:
        (exe_aluop_i == `MINIMIPS32_MFLO) ? lo_t: 
        (exe_aluop_i == `MINIMIPS32_MFC0) ? cp0_t:`ZERO_WORD;

   //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧妴luop闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳鐐
    assign arithres = 
        (exe_aluop_i == `MINIMIPS32_ADD  ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_LB   ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_LW   ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_SB   ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_SW   ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_SH   ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_ADDIU) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_SUBU ) ? (exe_src1_i + (~exe_src2_i) + 1):
        (exe_aluop_i == `MINIMIPS32_SLT  ) ? (($signed(exe_src1_i) < $signed(exe_src2_i)) ? 32'b1: 32'b0):
        (exe_aluop_i == `MINIMIPS32_ADDU ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_SUB  ) ? (exe_src1_i + (~exe_src2_i) + 1):
        (exe_aluop_i == `MINIMIPS32_SLTU ) ? (($unsigned(exe_src1_i) < $unsigned(exe_src2_i)) ? 32'b1 : 32'b0):
        (exe_aluop_i == `MINIMIPS32_ADDI ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_SLTI ) ? (($signed(exe_src1_i) < $signed(exe_src2_i)) ? 32'b1: 32'b0):
        (exe_aluop_i == `MINIMIPS32_SLTIU) ? ($unsigned(exe_src1_i) < $unsigned(exe_src2_i) ? 32'b1: 32'b0):
        (exe_aluop_i == `MINIMIPS32_LBU  ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_LH   ) ? (exe_src1_i + exe_src2_i):
        (exe_aluop_i == `MINIMIPS32_LHU  ) ? (exe_src1_i + exe_src2_i):`ZERO_WORD;
   //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧妴luop闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺屾稑鈻庡Ο杞扮暗缂備胶濮惧畷鐢靛垝閻㈠灚鍠嗛柛鏇ㄥ亽娴兼捇姊绘担鑺ョ《闁哥姵鍔欏鍛婄節濮橆剛顔嗛梺缁樺灱婵倝寮查幖浣圭厸闁稿本锚閳ь剚鐗滈埀顒佽壘缂嶅﹪寮婚妸鈺傚亜濠靛倸顦扮紞妤呮⒑閹稿海鈽夐柣顓炲€垮顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈崼鏇熲拺閻犳亽鍔岄弸鎴︽煛鐎ｎ亶鐓兼鐐茬箻閹藉酣宕掑⿰搴濈礃闂傚倷娴囧▔鏇㈠窗閺嶎灛鐔告媴閻戞ê顎涢柣鐔哥懃鐎氼剟顢旈敓锟�
    assign mulres           = ($signed(exe_src1_i) * $signed(exe_src2_i));
    assign mulures          =(exe_src1_i * exe_src2_i);

    assign exe_hilo_o = 
        (exe_aluop_i == `MINIMIPS32_MULTU)? mulures:
        (exe_aluop_i == `MINIMIPS32_MULT) ? mulres :
        (exe_aluop_i == `MINIMIPS32_DIV)  ? divres :
        (exe_aluop_i == `MINIMIPS32_DIVU)  ? divres :
        (exe_aluop_i == `MINIMIPS32_MTHI)  ? {exe_src1_i,exe_src1_i} :
        (exe_aluop_i == `MINIMIPS32_MTLO)  ? {exe_src1_i,exe_src1_i} : `ZERO_DWORD;

    assign exe_wa_o = exe_wa_i;
    assign exe_wreg_o = exe_wreg_i;



    //闂傚倷娴囧▔鏇㈠窗鎼淬們浜归柕濞у嫬顎涢柣鐔哥懃鐎氼剟顢旈崼鏇熲拺閻犳亽鍔岄弸娆愩亜椤愶綆娈滅€规洘鐟╂俊鍫曞幢濡ゅ﹣绱﹂梻鍌欐祰濞夋洟宕伴幇鏉垮嚑濠电姵鑹剧粻顖炴煟閹达絽袚闁哄懏鎮傞弻锟犲磼濡　鍋撻弽顐熷亾濮橆剛绉洪柡灞诲姂閹垽宕ㄦ繝鍕磿闂備礁缍婇ˉ鎾诲礂濮椻偓瀵偊骞樼拠鍙夘棟闂侀潧鐗嗗Λ妤咁敂閸洘鈷戦悹鎭掑妼閺嬫垿鏌＄€ｎ亶鐓兼鐐茬箻閹粓鎳為妷锔筋仧闂佽绻掗崑娑㈡晝閵堝鍋夐柨鐕傛嫹
    // wire [31:0] exe_src2_t =(exe_aluop_i==`MINIMIPS32_SUB)?(~exe_src2_i)+1 : exe_src2_i;
    // wire [31:0] arith_tmp=exe_src1_i+exe_src2_t;
    // wire [31:0] arith_tmp_2=exe_src1_i+exe_src2_i;
    // wire ov = (exe_aluop_i == `MINIMIPS32_SUB) ? ((!exe_src1_i[31] && !exe_src2_t[31] && arith_tmp[31]) || (exe_src1_i[31] && exe_src2_t[31] && !arith_tmp[31]))
    //            : (exe_aluop_i == `MINIMIPS32_ADD || exe_aluop_i == `MINIMIPS32_ADDI) ? 
    //            ((!exe_src1_i[31] && !exe_src2_i[31] && arith_tmp_2[31]) || (exe_src1_i[31] && exe_src2_i[31] && !arith_tmp_2[31])):0;
    
    wire ov = (exe_aluop_i == `MINIMIPS32_SUB) ? 
                   ((exe_src1_i[31] && !exe_src2_i[31] && !arithres[31])||(!exe_src1_i[31] && exe_src2_i[31] && arithres[31])) 
                   :
                   (exe_aluop_i == `MINIMIPS32_ADD || exe_aluop_i == `MINIMIPS32_ADDI) ? 
                       ((exe_src1_i[31] && exe_src2_i[31] && !arithres[31])||(!exe_src1_i[31] && !exe_src2_i[31] && arithres[31])) : 0;

    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш鐎殿噮鍓熼獮鍥嚋闂堟侗浼�
    assign exe_exccode_o =
        //(exe_aluop_i != `EXC_NONE) ? exe_exccode_i:
        ((exe_aluop_i==`MINIMIPS32_ADD|| exe_aluop_i==`MINIMIPS32_ADDI || exe_aluop_i==`MINIMIPS32_SUB)&&(ov==`TRUE_V))?`EXC_OV:exe_exccode_i;
    
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳槌栧妴lutype缂備胶铏庨崣搴ㄥ闯閿濆鏋侀柟鎹愵嚙濡﹢鏌曢崼婵囶棞妞ゅ繐鐖奸弻鐔虹箔濞戞ɑ澶勯柡鍛倐閺屾稑鈻庡Ο杞板枈濠碘槅鍨懗鍫曞箯鐎ｎ剚鍠嗛柛鏇ㄥ亽娴兼捇姊绘担鑺ョ《闁哥姵鍔欏鍛婄節濮橆剛顔嗛梺缁樺灱婵倝寮查崫銉х＜濠㈣泛锕ラ幉鍛娿亜閿濆骸娅嶆鐐茬箻閹粓鎳為妷锔筋仧闂備礁鎼崐鍫曞磹閺嶎偀鍋撳顒傜Ш闁哄被鍔戦幃銏ゅ川婵犲嫪绱曢梻浣哥秺椤ユ捇宕楀鈧顐﹀箻鐠囧弶顥濋梺闈涚墕濡顢旈敓锟�
    wire [2:0] alutype = exe_aluop_i[7:5];
    assign exe_wd_o = 
        (alutype == `MUL   ) ? mulres[31:0] : 
        (alutype == `LOGIC ) ? logicres :
        (alutype == `SHIFT ) ? shiftres :
        (alutype == `MOVE  ) ? moveres  :
        (alutype == `ARITH ) ? arithres : 
        (alutype == `JUMP  ) ? ret_addr : `ZERO_WORD;
    //闂傚倷娴囧▔鏇㈠窗閹版澘鍑犲┑鐘宠壘缁狀垶鏌ｉ幋锝呅撻柡鍛倐閺岋繝宕掑Ο琛″亾閺嶎偀鍋撳顒傜Ш鐎规洘绮岄鍏煎緞鐎ｎ偅顏熼梻浣告惈閸婂爼宕愰弽顐熷亾濮樼偓瀚�
    assign exe2id_wd = exe_wd_o;

endmodule